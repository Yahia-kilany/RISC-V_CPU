`timescale 1ns / 1ps

/*******************************************************************
*
* Module: inst_mem.v
* Project: RISC-V_CPU
* Author: Yahia Kilany
* Author: Ouail Slama 
* Description: 
*   Instruction memory module.
*   Provides 32-bit instructions for a 64-word memory.
*   Address input (addr_i) selects which instruction (data_o) to output asynchronous.
*
* Change history:
*   10/14/2025 – Initial lab version created
*   11/02/2025 – Adapted and cleaned for project use (Yahia)
*
*******************************************************************/

module inst_mem (
    input  wire [7:0]  addr_i, 
    output wire [31:0] data_o
);

    reg [31:0] mem_r [0:255];

    assign data_o = mem_r[addr_i];

    initial begin
mem_r[0]=32'b0000000_00000_00000_000_00000_0110011 ; //add x0, x0, x0
//added to be skipped since PC starts with 4 after reset
mem_r[1]=32'b000000000000_00000_010_00001_0000011 ; //lw x1, 0(x0)
mem_r[2]=32'b0000000_00000_00000_000_00000_0110011 ; //add x0, x0, x0
mem_r[3]=32'b0000000_00000_00000_000_00000_0110011 ; //add x0, x0, x0
mem_r[4]=32'b0000000_00000_00000_000_00000_0110011 ; //add x0, x0, x0
mem_r[5]=32'b000000000100_00000_010_00010_0000011 ; //lw x2, 4(x0)
mem_r[6]=32'b0000000_00000_00000_000_00000_0110011 ; //add x0, x0, x0
mem_r[7]=32'b0000000_00000_00000_000_00000_0110011 ; //add x0, x0, x0
mem_r[8]=32'b0000000_00000_00000_000_00000_0110011 ; //add x0, x0, x0
mem_r[9]=32'b000000001000_00000_010_00011_0000011 ; //lw x3, 8(x0)
mem_r[10]=32'b0000000_00000_00000_000_00000_0110011 ; //add x0, x0, x0
mem_r[11]=32'b0000000_00000_00000_000_00000_0110011 ; //add x0, x0, x0
mem_r[12]=32'b0000000_00000_00000_000_00000_0110011 ; //add x0, x0, x0
mem_r[13]=32'b0000000_00010_00001_110_00100_0110011 ; //or x4, x1, x2
mem_r[14]=32'b0000000_00000_00000_000_00000_0110011 ; //add x0, x0, x0
mem_r[15]=32'b0000000_00000_00000_000_00000_0110011 ; //add x0, x0, x0
mem_r[16]=32'b0000000_00000_00000_000_00000_0110011 ; //add x0, x0, x0
mem_r[17]=32'b0_000001_00011_00100_000_0000_0_1100011; //beq x4, x3, 16
mem_r[18]=32'b0000000_00000_00000_000_00000_0110011 ; //add x0, x0, x0
mem_r[19]=32'b0000000_00000_00000_000_00000_0110011 ; //add x0, x0, x0
mem_r[20]=32'b0000000_00000_00000_000_00000_0110011 ; //add x0, x0, x0
mem_r[21]=32'b0000000_00010_00001_000_00011_0110011 ; //add x3, x1, x2
mem_r[22]=32'b0000000_00000_00000_000_00000_0110011 ; //add x0, x0, x0
mem_r[23]=32'b0000000_00000_00000_000_00000_0110011 ; //add x0, x0, x0
mem_r[24]=32'b0000000_00000_00000_000_00000_0110011 ; //add x0, x0, x0
mem_r[25]=32'b0000000_00010_00011_000_00101_0110011 ; //add x5, x3, x2
mem_r[26]=32'b0000000_00000_00000_000_00000_0110011 ; //add x0, x0, x0
mem_r[27]=32'b0000000_00000_00000_000_00000_0110011 ; //add x0, x0, x0
mem_r[28]=32'b0000000_00000_00000_000_00000_0110011 ; //add x0, x0, x0
mem_r[29]=32'b0000000_00101_00000_010_01100_0100011; //sw x5, 12(x0)
mem_r[30]=32'b0000000_00000_00000_000_00000_0110011 ; //add x0, x0, x0
mem_r[31]=32'b0000000_00000_00000_000_00000_0110011 ; //add x0, x0, x0
mem_r[32]=32'b0000000_00000_00000_000_00000_0110011 ; //add x0, x0, x0
mem_r[33]=32'b000000001100_00000_010_00110_0000011 ; //lw x6, 12(x0)
mem_r[34]=32'b0000000_00000_00000_000_00000_0110011 ; //add x0, x0, x0
mem_r[35]=32'b0000000_00000_00000_000_00000_0110011 ; //add x0, x0, x0
mem_r[36]=32'b0000000_00000_00000_000_00000_0110011 ; //add x0, x0, x0
mem_r[37]=32'b0000000_00001_00110_111_00111_0110011 ; //and x7, x6, x1
mem_r[38]=32'b0000000_00000_00000_000_00000_0110011 ; //add x0, x0, x0
mem_r[39]=32'b0000000_00000_00000_000_00000_0110011 ; //add x0, x0, x0
mem_r[40]=32'b0000000_00000_00000_000_00000_0110011 ; //add x0, x0, x0
mem_r[41]=32'b0100000_00010_00001_000_01000_0110011 ; //sub x8, x1, x2
mem_r[42]=32'b0000000_00000_00000_000_00000_0110011 ; //add x0, x0, x0
mem_r[43]=32'b0000000_00000_00000_000_00000_0110011 ; //add x0, x0, x0
mem_r[44]=32'b0000000_00000_00000_000_00000_0110011 ; //add x0, x0, x0
mem_r[45]=32'b0000000_00010_00001_000_00000_0110011 ; //add x0, x1, x2
mem_r[46]=32'b0000000_00000_00000_000_00000_0110011 ; //add x0, x0, x0
mem_r[47]=32'b0000000_00000_00000_000_00000_0110011 ; //add x0, x0, x0
mem_r[48]=32'b0000000_00000_00000_000_00000_0110011 ; //add x0, x0, x0
mem_r[49]=32'b0000000_00001_00000_000_01001_0110011 ; //add x9, x0, x1    end

end 
endmodule